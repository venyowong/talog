module main

import core

pub struct TaggingLog {
pub mut:
	log string
	tags []core.Tag
}